module memoryStorage(
	input firstSign,
	input secondSign
	
);

endmodule 