module buttonDecode {
	input[3:0] KEY,
	input valid,
	input Clock_10ms,
	
	output backspace


};

always @ (posedge Clock_10ms)




